//**************************************************************************************************
// Project/Product : IDCT
// Description     : Inverse Discrete Cosine Transform 
//                   row and column 1D IDCT operation 
//                   with 3 stage pipeline in each 1D IDCT
// Dependencies    : global_defs.v, global_func.v, synch_fifo.v
// References      : 
//
//**************************************************************************************************
   
`timescale 1ns / 1ps

module add_en_12(
	clk_i,
	rst_n_i,

	data_1_i,
	data_2_i,
	data_sum_o,

	add_en_i,
	skip_neg_en_i
);


//----------------------------------------------------------------------------------------------------------------------
// Global constant and function headers
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// parameter definitions
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// localparam definitions
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// I/O signals
//----------------------------------------------------------------------------------------------------------------------

	// System Clock Signals
	input 															clk_i;
	input 															rst_n_i;

	input 				[11:0] 										data_1_i;
	input 				[11:0] 										data_2_i;
	output 	reg 		[11:0] 										data_sum_o;

	input 															add_en_i;
	input 															skip_neg_en_i;

//----------------------------------------------------------------------------------------------------------------------
// Internal wires and registers
//----------------------------------------------------------------------------------------------------------------------
			
	reg 				[11:0] 										r_add_1;
	reg 				[11:0] 										r_add_2;
	reg 				[11:0] 										r_add_3;
	reg 				[11:0] 										r_add_4;

	reg 															r_skip;

//----------------------------------------------------------------------------------------------------------------------
// Implmentation
//----------------------------------------------------------------------------------------------------------------------

	always @(posedge clk_i) begin 
		if(~rst_n_i) begin
			r_add_1 <= 0;
		end 
		else if(add_en_i) begin
			r_add_1[11:4] <= data_1_i[11:4] + data_2_i[11:4];
			r_add_1[3:0] <= 0;
		end
		else begin
			r_add_1 <= data_1_i;
		end
	end

	  always @(posedge clk_i) begin  : SKIP
	  	if(~rst_n_i) begin
	  		r_skip <= 0;
	  	end else begin
	  		r_skip <= skip_neg_en_i;
	  	end
	  end
//  
	  always @(posedge clk_i) begin : ADD_1
	  	if(~rst_n_i) begin
	  		r_add_2 <= 0;
	  	end 
	  	else if(r_skip && r_add_1[11:11] == 1) begin
	  		r_add_2 <= 0;
	  	end
	  	else begin
	  		r_add_2 <= r_add_1;
	  	end
	  end
//  
	  always @(posedge clk_i) begin : SUM
	  	if(~rst_n_i) begin
	  		r_add_3 <= 0;
	  		r_add_4 <= 0;
	  		data_sum_o <= 0;
	  	end 
	  	else begin
	  		r_add_3 <= r_add_2;
	  		r_add_4 <= r_add_3;
	  		data_sum_o <= r_add_4;
	  	end
	  end

//----------------------------------------------------------------------------------------------------------------------
// Sub module instantiation
//----------------------------------------------------------------------------------------------------------------------

	
endmodule

