//**************************************************************************************************
// Project/Product : IDCT
// Description     : Inverse Discrete Cosine Transform 
//                   row and column 1D IDCT operation 
//                   with 3 stage pipeline in each 1D IDCT
// Dependencies    : global_defs.v, global_func.v, synch_fifo.v
// References      : 
//
//**************************************************************************************************
   
`timescale 1ns / 1ps

module expand_add(
	clk_i,
	rst_n_i,

	expand_1_i,
	expand_2_i,
	expand_sum_o,

	add_en_i
);


//----------------------------------------------------------------------------------------------------------------------
// Global constant and function headers
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// parameter definitions
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// localparam definitions
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// I/O signals
//----------------------------------------------------------------------------------------------------------------------

	// System Clock Signals
	input 															clk_i;
	input 															rst_n_i;

	// Add control Signals
	input 					[47:0] 									expand_1_i;
	input 					[47:0] 									expand_2_i;
	output 					[47:0] 									expand_sum_o;

	input 															add_en_i;

//----------------------------------------------------------------------------------------------------------------------
// Internal wires and registers
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// Implmentation
//----------------------------------------------------------------------------------------------------------------------

//----------------------------------------------------------------------------------------------------------------------
// Sub module instantiation
//----------------------------------------------------------------------------------------------------------------------

	add_en_12 float_add_1_inst
	(
		.clk_i 								(clk_i),
		.rst_n_i 							(rst_n_i),

		.data_1_i 							(expand_1_i[47:36]),
		.data_2_i 							(expand_2_i[47:36]),
		.data_sum_o 						(expand_sum_o[47:36]),

		.add_en_i 							(add_en_i),
		.skip_neg_en_i 						(0)
	);

	// Float ADD 2 Instantiation
	add_en_12 float_add_2_inst
	(
		.clk_i 				 				(clk_i),
		.rst_n_i 							(rst_n_i),

		.data_1_i 							(expand_1_i[35:24]),
		.data_2_i 							(expand_2_i[35:24]),
		.data_sum_o 						(expand_sum_o[35:24]),

		.add_en_i 							(add_en_i),
		.skip_neg_en_i 						(0)
	);

	// Float ADD 3 Instantiation
	add_en_12 float_add_3_inst
	(
		.clk_i 				 				(clk_i),
		.rst_n_i 							(rst_n_i),

		.data_1_i 							(expand_1_i[23:12]),
		.data_2_i 							(expand_2_i[23:12]),
		.data_sum_o 						(expand_sum_o[23:12]),

		.add_en_i 							(add_en_i),
		.skip_neg_en_i 						(0)
	);

	// Float ADD 4 Instantiation
	add_en_12 float_add_4_inst
	(
		.clk_i 				 				(clk_i),
		.rst_n_i 							(rst_n_i),

		.data_1_i 							(expand_1_i[11:00]),
		.data_2_i 							(expand_2_i[11:00]),
		.data_sum_o 						(expand_sum_o[11:00]),

		.add_en_i 							(add_en_i),
		.skip_neg_en_i 						(0)
	);

endmodule

